library ieee;
use ieee.std_logic_1164.all;

entity abcExpr_tb_CU is
    port (
        reset_n,
        clock,
        start: in std_logic;
        
    );